// Copyright (c) 2024 Princeton University
// All rights reserved.
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//     * Redistributions of source code must retain the above copyright
//       notice, this list of conditions and the following disclaimer.
//     * Redistributions in binary form must reproduce the above copyright
//       notice, this list of conditions and the following disclaimer in the
//       documentation and/or other materials provided with the distribution.
//     * Neither the name of the copyright holder nor the
//       names of its contributors may be used to endorse or promote products
//       derived from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.


// Automatically generated by PRGA's RTL generator
`ifndef PRGA_PKTCHAIN_SYSTEM_H
`define PRGA_PKTCHAIN_SYSTEM_H

`include "prga_system.vh"
`include "pktchain.vh"

`define PRGA_CREG_ADDR_PKTCHAIN_BITSTREAM_FIFO      `PRGA_CREG_ADDR_WIDTH'h900  //  64b

`define PRGA_EFLAGS_PKTCHAIN_RESP_INVAL             32
`define PRGA_EFLAGS_PKTCHAIN_BITSTREAM_CORRUPTED    33
`define PRGA_EFLAGS_PKTCHAIN_BITSTREAM_INCOMPLETE   34
`define PRGA_EFLAGS_PKTCHAIN_BITSTREAM_REDUNDANT    35

`endif /* PRGA_PKTCHAIN_SYSTEM_H */